`timescale 1ns / 1ps

module half_adder_structural(sum,carry,a,b);
output sum,carry;
input a,b;

xor s(sum,a,b);
and cout(carry,a,b);
endmodule
